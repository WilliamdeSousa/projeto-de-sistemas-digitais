// exemplo dado por George em aula remota

module hello();
  initial begin
    $display("*** Hello World ***");
    $finish();
  end
endmodule: hello;